module FD_Testbench ();

endmodule 